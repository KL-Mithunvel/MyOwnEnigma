`timescale 1ns / 1ps
//module blinky(
//    input clk,
//    output led,
//    input sw
//    );
//    reg [24:0] count = 0;  
//    assign led = count[24];
//    always @ (posedge(clk)) count <= count + 1;
//endmodule
